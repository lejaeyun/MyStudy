module RippleCarryAdder_tb;

reg A0;
reg A1;
reg A2;
reg A3;
reg B0;
reg B1;
reg B2;
reg B3;
reg C0;
wire C4;
wire S0;
wire S1;
wire S2;
wire S3;

Ripple_Carry_Adder
 U0 (
  .A0(A0),
  .A1(A1),
  .A2(A2),
  .A3(A3),
  .B0(B0),
  .B1(B1),
  .B2(B2),
  .B3(B3),
  .C0(C0),
  .C4(C4),
  .S0(S0),
  .S1(S1),
  .S2(S2),
  .S3(S3));

  initial
  begin
    A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b0;
    #100 A0 = 1'b1;
    #100 A0 = 1'b0;

  end

  initial
  begin
    A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;
    #100 A1 = 1'b1;
    #100 A1 = 1'b0;

  end

  initial
  begin
    A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;
    #100 A2 = 1'b1;
    #100 A2 = 1'b0;

  end

  initial
  begin
    A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;
    #100 A3 = 1'b1;
    #100 A3 = 1'b0;

  end

  initial
  begin
    B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;
    #100 B0 = 1'b1;
    #100 B0 = 1'b0;

  end

  initial
  begin
    B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;
    #100 B1 = 1'b1;
    #100 B1 = 1'b0;

  end

  initial
  begin
    B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;
    #100 B2 = 1'b1;
    #100 B2 = 1'b0;

  end

  initial
  begin
    B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;
    #100 B3 = 1'b1;
    #100 B3 = 1'b0;

  end

  initial
  begin
    C0 = 1'b0;
  end

endmodule
